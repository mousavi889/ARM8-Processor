module reg_bank(clk, rst, raddr1, raddr2, waddr, din, dout1, dout2, regwrite);
	input 			clk;
	input 			rst;
	input 	[4:0] 	raddr1;
	input 	[4:0] 	raddr2;
	input 	[4:0] 	waddr;
	input 			regwrite;
	input 	[31:0] 	din;
	output 	[31:0] 	dout1;
	reg    	[31:0] 	dout1;
	output 	[31:0] 	dout2;
	reg    	[31:0] 	dout2;
	reg    	[31:0] 	bank [0:31];
	always @(raddr1)
		dout1 = bank[raddr1];
	always @(raddr2)
		dout2 = bank[raddr2];
    always @ (rst or posedge clk)
    begin
      if (rst)
			begin
				bank[0] = 32'b00000000000000000000000000000001;
				bank[1] = 32'b00000000000000000000000000000011;
				bank[2] = 32'b00000000000000000000000000000000;
				bank[3] = 32'b00000000000000000000000000000000;
				bank[4] = 32'b00000000000000000000000000000000;
				bank[5] = 32'b00000000000000000000000000000000;
				bank[6] = 32'b00000000000000000000000000000000;
				bank[7] = 32'b00000000000000000000000000000000;
				bank[8] = 32'b00000000000000000000000000000000;
				bank[9] = 32'b00000000000000000000000000000000;
				bank[10] = 32'b00000000000000000000000000000000;
				bank[11] = 32'b00000000000000000000000000000000;
				bank[12] = 32'b00000000000000000000000000000000;
				bank[13] = 32'b00000000000000000000000000000000;
				bank[14] = 32'b00000000000000000000000000000000;
				bank[15] = 32'b00000000000000000000000000000000;
				bank[16] = 32'b00000000000000000000000000000000;
				bank[17] = 32'b00000000000000000000000000000000;
				bank[18] = 32'b00000000000000000000000000000000;
				bank[19] = 32'b00000000000000000000000000000000;
				bank[20] = 32'b00000000000000000000000000000000;
				bank[21] = 32'b00000000000000000000000000000000;
				bank[22] = 32'b00000000000000000000000000000000;
				bank[23] = 32'b00000000000000000000000000000000;
				bank[24] = 32'b00000000000000000000000000000000;
				bank[25] = 32'b00000000000000000000000000000000;
				bank[26] = 32'b00000000000000000000000000000000;
				bank[27] = 32'b00000000000000000000000000000000;
				bank[28] = 32'b00000000000000000000000000000000;
				bank[29] = 32'b00000000000000000000000000000000;
				bank[30] = 32'b00000000000000000000000000000000;
				bank[31] = 32'b00000000000000000000000000000000;
			end
      else if (clk)
			if (regwrite)
				bank[waddr] = din;
	end
endmodule
